library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.all;
USE work.LED_matrix_type_package.ALL;

entity TestPattern is
    Port ( clk : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           addr_out : out  STD_LOGIC_VECTOR (3 downto 0);
           oe : out  STD_LOGIC;
           latch : out  STD_LOGIC;
           r0 : out  STD_LOGIC;
           g0 : out  STD_LOGIC;
           b0 : out  STD_LOGIC;
           r1 : out  STD_LOGIC;
           g1 : out  STD_LOGIC;
           b1 : out  STD_LOGIC;
           sclk : out  STD_LOGIC);
end TestPattern;

architecture Behavioral of TestPattern is

	COMPONENT LEDMatrixDriver
	PORT(
		clk : IN std_logic;
		data : IN RGB_LED_array;
		rst : IN std_logic;     
		pwm_mode : in  STD_LOGIC;		
		sclk : OUT std_logic;
		r0 : OUT std_logic;
		g0 : OUT std_logic;
		b0 : OUT std_logic;
		r1 : OUT std_logic;
		g1 : OUT std_logic;
		b1 : OUT std_logic;
		oe : OUT std_logic;
		latch : OUT std_logic;
		addr_out : OUT std_logic_vector(3 downto 0)
		);
	END COMPONENT;
	
	signal data0: RGB_LED_array;
	
	signal counter: unsigned(4 downto 0);
	signal counter2: unsigned(4 downto 0);
	
begin

				data0(0) <= (
					( "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000" ),
					( "00000000", "00000000", "00000000", "00000000", "00000000", "00000001", "00000001", "00000001", "00000001", "00000010", "00000010", "00000010", "00000010", "00000011", "00000011", "00000011", "00000011", "00000100", "00000100", "00000100", "00000100", "00000101", "00000101", "00000101", "00000101", "00000110", "00000110", "00000110", "00000110", "00000111", "00000111", "00000111" ),
					( "00000000", "00000000", "00000000", "00000001", "00000001", "00000010", "00000010", "00000011", "00000011", "00000100", "00000100", "00000101", "00000101", "00000110", "00000110", "00000111", "00000111", "00001000", "00001000", "00001001", "00001001", "00001010", "00001010", "00001011", "00001011", "00001100", "00001100", "00001101", "00001101", "00001110", "00001110", "00001111" ),
					( "00000000", "00000000", "00000001", "00000010", "00000010", "00000011", "00000100", "00000101", "00000101", "00000110", "00000111", "00001000", "00001000", "00001001", "00001010", "00001011", "00001011", "00001100", "00001101", "00001110", "00001110", "00001111", "00010000", "00010001", "00010001", "00010010", "00010011", "00010100", "00010100", "00010101", "00010110", "00010111" ),
					( "00000000", "00000000", "00000001", "00000010", "00000011", "00000100", "00000101", "00000110", "00000111", "00001000", "00001001", "00001010", "00001011", "00001100", "00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", "00011101", "00011110" ),
					( "00000000", "00000001", "00000010", "00000011", "00000100", "00000110", "00000111", "00001000", "00001001", "00001011", "00001100", "00001101", "00001110", "00010000", "00010001", "00010010", "00010011", "00010101", "00010110", "00010111", "00011000", "00011010", "00011011", "00011100", "00011101", "00011111", "00100000", "00100001", "00100010", "00100100", "00100101", "00100110" ),
					( "00000000", "00000001", "00000010", "00000100", "00000101", "00000111", "00001000", "00001010", "00001011", "00001101", "00001110", "00010000", "00010001", "00010011", "00010100", "00010110", "00010111", "00011001", "00011010", "00011100", "00011101", "00011111", "00100000", "00100010", "00100011", "00100101", "00100110", "00101000", "00101001", "00101011", "00101100", "00101110" ),
					( "00000000", "00000001", "00000011", "00000101", "00000110", "00001000", "00001010", "00001100", "00001101", "00001111", "00010001", "00010011", "00010100", "00010110", "00011000", "00011010", "00011011", "00011101", "00011111", "00100001", "00100010", "00100100", "00100110", "00101000", "00101001", "00101011", "00101101", "00101111", "00110000", "00110010", "00110100", "00110110" ),
					( "00000000", "00000001", "00000011", "00000101", "00000111", "00001001", "00001011", "00001101", "00001111", "00010001", "00010011", "00010101", "00010111", "00011001", "00011011", "00011101", "00011111", "00100001", "00100011", "00100101", "00100111", "00101001", "00101011", "00101101", "00101111", "00110001", "00110011", "00110101", "00110111", "00111001", "00111011", "00111101" ),
					( "00000000", "00000010", "00000100", "00000110", "00001000", "00001011", "00001101", "00001111", "00010001", "00010100", "00010110", "00011000", "00011010", "00011101", "00011111", "00100001", "00100011", "00100110", "00101000", "00101010", "00101100", "00101111", "00110001", "00110011", "00110101", "00111000", "00111010", "00111100", "00111110", "01000000", "01000011", "01000101" ),
					( "00000000", "00000010", "00000100", "00000111", "00001001", "00001100", "00001110", "00010001", "00010011", "00010110", "00011000", "00011011", "00011101", "00100000", "00100010", "00100101", "00100111", "00101010", "00101100", "00101111", "00110001", "00110100", "00110110", "00111001", "00111011", "00111110", "01000000", "01000011", "01000101", "01001000", "01001010", "01001101" ),
					( "00000000", "00000010", "00000101", "00001000", "00001010", "00001101", "00010000", "00010011", "00010101", "00011000", "00011011", "00011110", "00100000", "00100011", "00100110", "00101001", "00101011", "00101110", "00110001", "00110100", "00110110", "00111001", "00111100", "00111111", "01000001", "01000100", "01000111", "01001001", "01001100", "01001111", "01010010", "01010100" ),
					( "00000000", "00000010", "00000101", "00001000", "00001011", "00001110", "00010001", "00010100", "00010111", "00011010", "00011101", "00100000", "00100011", "00100110", "00101001", "00101100", "00101111", "00110010", "00110101", "00111000", "00111011", "00111110", "01000001", "01000100", "01000111", "01001010", "01001101", "01010000", "01010011", "01010110", "01011001", "01011100" ),
					( "00000000", "00000011", "00000110", "00001001", "00001100", "00010000", "00010011", "00010110", "00011001", "00011101", "00100000", "00100011", "00100110", "00101010", "00101101", "00110000", "00110011", "00110111", "00111010", "00111101", "01000000", "01000011", "01000111", "01001010", "01001101", "01010000", "01010100", "01010111", "01011010", "01011101", "01100001", "01100100" ),
					( "00000000", "00000011", "00000110", "00001010", "00001101", "00010001", "00010100", "00011000", "00011011", "00011111", "00100010", "00100110", "00101001", "00101101", "00110000", "00110100", "00110111", "00111011", "00111110", "01000010", "01000101", "01001001", "01001100", "01010000", "01010011", "01010111", "01011010", "01011110", "01100001", "01100101", "01101000", "01101100" ),
					( "00000000", "00000011", "00000111", "00001011", "00001110", "00010010", "00010110", "00011010", "00011101", "00100001", "00100101", "00101001", "00101100", "00110000", "00110100", "00111000", "00111011", "00111111", "01000011", "01000110", "01001010", "01001110", "01010010", "01010101", "01011001", "01011101", "01100001", "01100100", "01101000", "01101100", "01110000", "01110011" ),
					( "00000000", "00000011", "00000111", "00001011", "00001111", "00010011", "00010111", "00011011", "00011111", "00100011", "00100111", "00101011", "00101111", "00110011", "00110111", "00111011", "00111111", "01000011", "01000111", "01001011", "01001111", "01010011", "01010111", "01011011", "01011111", "01100011", "01100111", "01101011", "01101111", "01110011", "01110111", "01111011" ),
					( "00000000", "00000100", "00001000", "00001100", "00010000", "00010101", "00011001", "00011101", "00100001", "00100110", "00101010", "00101110", "00110010", "00110111", "00111011", "00111111", "01000011", "01000111", "01001100", "01010000", "01010100", "01011000", "01011101", "01100001", "01100101", "01101001", "01101110", "01110010", "01110110", "01111010", "01111111", "10000011" ),
					( "00000000", "00000100", "00001000", "00001101", "00010001", "00010110", "00011010", "00011111", "00100011", "00101000", "00101100", "00110001", "00110101", "00111010", "00111110", "01000011", "01000111", "01001100", "01010000", "01010101", "01011001", "01011110", "01100010", "01100111", "01101011", "01110000", "01110100", "01111001", "01111101", "10000001", "10000110", "10001010" ),
					( "00000000", "00000100", "00001001", "00001110", "00010010", "00010111", "00011100", "00100001", "00100101", "00101010", "00101111", "00110100", "00111000", "00111101", "01000010", "01000110", "01001011", "01010000", "01010101", "01011001", "01011110", "01100011", "01101000", "01101100", "01110001", "01110110", "01111011", "01111111", "10000100", "10001001", "10001101", "10010010" ),
					( "00000000", "00000100", "00001001", "00001110", "00010011", "00011000", "00011101", "00100010", "00100111", "00101100", "00110001", "00110110", "00111011", "01000000", "01000101", "01001010", "01001111", "01010100", "01011001", "01011110", "01100011", "01101000", "01101101", "01110010", "01110111", "01111100", "10000001", "10000110", "10001011", "10010000", "10010101", "10011010" ),
					( "00000000", "00000101", "00001010", "00001111", "00010100", "00011010", "00011111", "00100100", "00101001", "00101111", "00110100", "00111001", "00111110", "01000011", "01001001", "01001110", "01010011", "01011000", "01011110", "01100011", "01101000", "01101101", "01110011", "01111000", "01111101", "10000010", "10000111", "10001101", "10010010", "10010111", "10011100", "10100010" ),
					( "00000000", "00000101", "00001010", "00010000", "00010101", "00011011", "00100000", "00100110", "00101011", "00110001", "00110110", "00111100", "01000001", "01000111", "01001100", "01010010", "01010111", "01011101", "01100010", "01101000", "01101101", "01110011", "01111000", "01111110", "10000011", "10001000", "10001110", "10010011", "10011001", "10011110", "10100100", "10101001" ),
					( "00000000", "00000101", "00001011", "00010001", "00010110", "00011100", "00100010", "00101000", "00101101", "00110011", "00111001", "00111111", "01000100", "01001010", "01010000", "01010101", "01011011", "01100001", "01100111", "01101100", "01110010", "01111000", "01111110", "10000011", "10001001", "10001111", "10010100", "10011010", "10100000", "10100110", "10101011", "10110001" ),
					( "00000000", "00000101", "00001011", "00010001", "00010111", "00011101", "00100011", "00101001", "00101111", "00110101", "00111011", "01000001", "01000111", "01001101", "01010011", "01011001", "01011111", "01100101", "01101011", "01110001", "01110111", "01111101", "10000011", "10001001", "10001111", "10010101", "10011011", "10100001", "10100111", "10101101", "10110011", "10111001" ),
					( "00000000", "00000110", "00001100", "00010010", "00011000", "00011111", "00100101", "00101011", "00110001", "00111000", "00111110", "01000100", "01001010", "01010000", "01010111", "01011101", "01100011", "01101001", "01110000", "01110110", "01111100", "10000010", "10001000", "10001111", "10010101", "10011011", "10100001", "10101000", "10101110", "10110100", "10111010", "11000000" ),
					( "00000000", "00000110", "00001100", "00010011", "00011001", "00100000", "00100110", "00101101", "00110011", "00111010", "01000000", "01000111", "01001101", "01010100", "01011010", "01100001", "01100111", "01101110", "01110100", "01111011", "10000001", "10000111", "10001110", "10010100", "10011011", "10100001", "10101000", "10101110", "10110101", "10111011", "11000010", "11001000" ),
					( "00000000", "00000110", "00001101", "00010100", "00011010", "00100001", "00101000", "00101111", "00110101", "00111100", "01000011", "01001001", "01010000", "01010111", "01011110", "01100100", "01101011", "01110010", "01111001", "01111111", "10000110", "10001101", "10010011", "10011010", "10100001", "10101000", "10101110", "10110101", "10111100", "11000010", "11001001", "11010000" ),
					( "00000000", "00000110", "00001101", "00010100", "00011011", "00100010", "00101001", "00110000", "00110111", "00111110", "01000101", "01001100", "01010011", "01011010", "01100001", "01101000", "01101111", "01110110", "01111101", "10000100", "10001011", "10010010", "10011001", "10100000", "10100111", "10101110", "10110101", "10111100", "11000011", "11001010", "11010001", "11011000" ),
					( "00000000", "00000111", "00001110", "00010101", "00011100", "00100100", "00101011", "00110010", "00111001", "01000000", "01001000", "01001111", "01010110", "01011101", "01100101", "01101100", "01110011", "01111010", "10000001", "10001001", "10010000", "10010111", "10011110", "10100110", "10101101", "10110100", "10111011", "11000010", "11001010", "11010001", "11011000", "11011111" ),
					( "00000000", "00000111", "00001110", "00010110", "00011101", "00100101", "00101100", "00110100", "00111011", "01000011", "01001010", "01010010", "01011001", "01100001", "01101000", "01110000", "01110111", "01111111", "10000110", "10001101", "10010101", "10011100", "10100100", "10101011", "10110011", "10111010", "11000010", "11001001", "11010001", "11011000", "11100000", "11100111" ),
					( "00000000", "00000111", "00001111", "00010111", "00011110", "00100110", "00101110", "00110110", "00111101", "01000101", "01001101", "01010100", "01011100", "01100100", "01101100", "01110011", "01111011", "10000011", "10001010", "10010010", "10011010", "10100010", "10101001", "10110001", "10111001", "11000000", "11001000", "11010000", "11011000", "11011111", "11100111", "11101111" )
				);
					
				data0(1) <= (
					( "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000" ),
					( "00000111", "00000111", "00000111", "00000110", "00000110", "00000110", "00000110", "00000101", "00000101", "00000101", "00000101", "00000100", "00000100", "00000100", "00000100", "00000011", "00000011", "00000011", "00000011", "00000010", "00000010", "00000010", "00000010", "00000001", "00000001", "00000001", "00000001", "00000000", "00000000", "00000000", "00000000", "00000000" ),
					( "00001111", "00001110", "00001110", "00001101", "00001101", "00001100", "00001100", "00001011", "00001011", "00001010", "00001010", "00001001", "00001001", "00001000", "00001000", "00000111", "00000111", "00000110", "00000110", "00000101", "00000101", "00000100", "00000100", "00000011", "00000011", "00000010", "00000010", "00000001", "00000001", "00000000", "00000000", "00000000" ),
					( "00010111", "00010110", "00010101", "00010100", "00010100", "00010011", "00010010", "00010001", "00010001", "00010000", "00001111", "00001110", "00001110", "00001101", "00001100", "00001011", "00001011", "00001010", "00001001", "00001000", "00001000", "00000111", "00000110", "00000101", "00000101", "00000100", "00000011", "00000010", "00000010", "00000001", "00000000", "00000000" ),
					( "00011110", "00011101", "00011100", "00011011", "00011010", "00011001", "00011000", "00010111", "00010110", "00010101", "00010100", "00010011", "00010010", "00010001", "00010000", "00001111", "00001110", "00001101", "00001100", "00001011", "00001010", "00001001", "00001000", "00000111", "00000110", "00000101", "00000100", "00000011", "00000010", "00000001", "00000000", "00000000" ),
					( "00100110", "00100101", "00100100", "00100010", "00100001", "00100000", "00011111", "00011101", "00011100", "00011011", "00011010", "00011000", "00010111", "00010110", "00010101", "00010011", "00010010", "00010001", "00010000", "00001110", "00001101", "00001100", "00001011", "00001001", "00001000", "00000111", "00000110", "00000100", "00000011", "00000010", "00000001", "00000000" ),
					( "00101110", "00101100", "00101011", "00101001", "00101000", "00100110", "00100101", "00100011", "00100010", "00100000", "00011111", "00011101", "00011100", "00011010", "00011001", "00010111", "00010110", "00010100", "00010011", "00010001", "00010000", "00001110", "00001101", "00001011", "00001010", "00001000", "00000111", "00000101", "00000100", "00000010", "00000001", "00000000" ),
					( "00110110", "00110100", "00110010", "00110000", "00101111", "00101101", "00101011", "00101001", "00101000", "00100110", "00100100", "00100010", "00100001", "00011111", "00011101", "00011011", "00011010", "00011000", "00010110", "00010100", "00010011", "00010001", "00001111", "00001101", "00001100", "00001010", "00001000", "00000110", "00000101", "00000011", "00000001", "00000000" ),
					( "00111101", "00111011", "00111001", "00110111", "00110101", "00110011", "00110001", "00101111", "00101101", "00101011", "00101001", "00100111", "00100101", "00100011", "00100001", "00011111", "00011101", "00011011", "00011001", "00010111", "00010101", "00010011", "00010001", "00001111", "00001101", "00001011", "00001001", "00000111", "00000101", "00000011", "00000001", "00000000" ),
					( "01000101", "01000011", "01000000", "00111110", "00111100", "00111010", "00111000", "00110101", "00110011", "00110001", "00101111", "00101100", "00101010", "00101000", "00100110", "00100011", "00100001", "00011111", "00011101", "00011010", "00011000", "00010110", "00010100", "00010001", "00001111", "00001101", "00001011", "00001000", "00000110", "00000100", "00000010", "00000000" ),
					( "01001101", "01001010", "01001000", "01000101", "01000011", "01000000", "00111110", "00111011", "00111001", "00110110", "00110100", "00110001", "00101111", "00101100", "00101010", "00100111", "00100101", "00100010", "00100000", "00011101", "00011011", "00011000", "00010110", "00010011", "00010001", "00001110", "00001100", "00001001", "00000111", "00000100", "00000010", "00000000" ),
					( "01010100", "01010010", "01001111", "01001100", "01001001", "01000111", "01000100", "01000001", "00111111", "00111100", "00111001", "00110110", "00110100", "00110001", "00101110", "00101011", "00101001", "00100110", "00100011", "00100000", "00011110", "00011011", "00011000", "00010101", "00010011", "00010000", "00001101", "00001010", "00001000", "00000101", "00000010", "00000000" ),
					( "01011100", "01011001", "01010110", "01010011", "01010000", "01001101", "01001010", "01000111", "01000100", "01000001", "00111110", "00111011", "00111000", "00110101", "00110010", "00101111", "00101100", "00101001", "00100110", "00100011", "00100000", "00011101", "00011010", "00010111", "00010100", "00010001", "00001110", "00001011", "00001000", "00000101", "00000010", "00000000" ),
					( "01100100", "01100001", "01011101", "01011010", "01010111", "01010100", "01010000", "01001101", "01001010", "01000111", "01000011", "01000000", "00111101", "00111010", "00110111", "00110011", "00110000", "00101101", "00101010", "00100110", "00100011", "00100000", "00011101", "00011001", "00010110", "00010011", "00010000", "00001100", "00001001", "00000110", "00000011", "00000000" ),
					( "01101100", "01101000", "01100101", "01100001", "01011110", "01011010", "01010111", "01010011", "01010000", "01001100", "01001001", "01000101", "01000010", "00111110", "00111011", "00110111", "00110100", "00110000", "00101101", "00101001", "00100110", "00100010", "00011111", "00011011", "00011000", "00010100", "00010001", "00001101", "00001010", "00000110", "00000011", "00000000" ),
					( "01110011", "01110000", "01101100", "01101000", "01100100", "01100001", "01011101", "01011001", "01010101", "01010010", "01001110", "01001010", "01000110", "01000011", "00111111", "00111011", "00111000", "00110100", "00110000", "00101100", "00101001", "00100101", "00100001", "00011101", "00011010", "00010110", "00010010", "00001110", "00001011", "00000111", "00000011", "00000000" ),
					( "01111011", "01110111", "01110011", "01101111", "01101011", "01100111", "01100011", "01011111", "01011011", "01010111", "01010011", "01001111", "01001011", "01000111", "01000011", "00111111", "00111011", "00110111", "00110011", "00101111", "00101011", "00100111", "00100011", "00011111", "00011011", "00010111", "00010011", "00001111", "00001011", "00000111", "00000011", "00000000" ),
					( "10000011", "01111111", "01111010", "01110110", "01110010", "01101110", "01101001", "01100101", "01100001", "01011101", "01011000", "01010100", "01010000", "01001100", "01000111", "01000011", "00111111", "00111011", "00110111", "00110010", "00101110", "00101010", "00100110", "00100001", "00011101", "00011001", "00010101", "00010000", "00001100", "00001000", "00000100", "00000000" ),
					( "10001010", "10000110", "10000001", "01111101", "01111001", "01110100", "01110000", "01101011", "01100111", "01100010", "01011110", "01011001", "01010101", "01010000", "01001100", "01000111", "01000011", "00111110", "00111010", "00110101", "00110001", "00101100", "00101000", "00100011", "00011111", "00011010", "00010110", "00010001", "00001101", "00001000", "00000100", "00000000" ),
					( "10010010", "10001101", "10001001", "10000100", "01111111", "01111011", "01110110", "01110001", "01101100", "01101000", "01100011", "01011110", "01011001", "01010101", "01010000", "01001011", "01000110", "01000010", "00111101", "00111000", "00110100", "00101111", "00101010", "00100101", "00100001", "00011100", "00010111", "00010010", "00001110", "00001001", "00000100", "00000000" ),
					( "10011010", "10010101", "10010000", "10001011", "10000110", "10000001", "01111100", "01110111", "01110010", "01101101", "01101000", "01100011", "01011110", "01011001", "01010100", "01001111", "01001010", "01000101", "01000000", "00111011", "00110110", "00110001", "00101100", "00100111", "00100010", "00011101", "00011000", "00010011", "00001110", "00001001", "00000100", "00000000" ),
					( "10100010", "10011100", "10010111", "10010010", "10001101", "10000111", "10000010", "01111101", "01111000", "01110011", "01101101", "01101000", "01100011", "01011110", "01011000", "01010011", "01001110", "01001001", "01000011", "00111110", "00111001", "00110100", "00101111", "00101001", "00100100", "00011111", "00011010", "00010100", "00001111", "00001010", "00000101", "00000000" ),
					( "10101001", "10100100", "10011110", "10011001", "10010011", "10001110", "10001000", "10000011", "01111110", "01111000", "01110011", "01101101", "01101000", "01100010", "01011101", "01010111", "01010010", "01001100", "01000111", "01000001", "00111100", "00110110", "00110001", "00101011", "00100110", "00100000", "00011011", "00010101", "00010000", "00001010", "00000101", "00000000" ),
					( "10110001", "10101011", "10100110", "10100000", "10011010", "10010100", "10001111", "10001001", "10000011", "01111110", "01111000", "01110010", "01101100", "01100111", "01100001", "01011011", "01010101", "01010000", "01001010", "01000100", "00111111", "00111001", "00110011", "00101101", "00101000", "00100010", "00011100", "00010110", "00010001", "00001011", "00000101", "00000000" ),
					( "10111001", "10110011", "10101101", "10100111", "10100001", "10011011", "10010101", "10001111", "10001001", "10000011", "01111101", "01110111", "01110001", "01101011", "01100101", "01011111", "01011001", "01010011", "01001101", "01000111", "01000001", "00111011", "00110101", "00101111", "00101001", "00100011", "00011101", "00010111", "00010001", "00001011", "00000101", "00000000" ),
					( "11000000", "10111010", "10110100", "10101110", "10101000", "10100001", "10011011", "10010101", "10001111", "10001000", "10000010", "01111100", "01110110", "01110000", "01101001", "01100011", "01011101", "01010111", "01010000", "01001010", "01000100", "00111110", "00111000", "00110001", "00101011", "00100101", "00011111", "00011000", "00010010", "00001100", "00000110", "00000000" ),
					( "11001000", "11000010", "10111011", "10110101", "10101110", "10101000", "10100001", "10011011", "10010100", "10001110", "10000111", "10000001", "01111011", "01110100", "01101110", "01100111", "01100001", "01011010", "01010100", "01001101", "01000111", "01000000", "00111010", "00110011", "00101101", "00100110", "00100000", "00011001", "00010011", "00001100", "00000110", "00000000" ),
					( "11010000", "11001001", "11000010", "10111100", "10110101", "10101110", "10101000", "10100001", "10011010", "10010011", "10001101", "10000110", "01111111", "01111001", "01110010", "01101011", "01100100", "01011110", "01010111", "01010000", "01001001", "01000011", "00111100", "00110101", "00101111", "00101000", "00100001", "00011010", "00010100", "00001101", "00000110", "00000000" ),
					( "11011000", "11010001", "11001010", "11000011", "10111100", "10110101", "10101110", "10100111", "10100000", "10011001", "10010010", "10001011", "10000100", "01111101", "01110110", "01101111", "01101000", "01100001", "01011010", "01010011", "01001100", "01000101", "00111110", "00110111", "00110000", "00101001", "00100010", "00011011", "00010100", "00001101", "00000110", "00000000" ),
					( "11011111", "11011000", "11010001", "11001010", "11000010", "10111011", "10110100", "10101101", "10100110", "10011110", "10010111", "10010000", "10001001", "10000001", "01111010", "01110011", "01101100", "01100101", "01011101", "01010110", "01001111", "01001000", "01000000", "00111001", "00110010", "00101011", "00100100", "00011100", "00010101", "00001110", "00000111", "00000000" ),
					( "11100111", "11100000", "11011000", "11010001", "11001001", "11000010", "10111010", "10110011", "10101011", "10100100", "10011100", "10010101", "10001101", "10000110", "01111111", "01110111", "01110000", "01101000", "01100001", "01011001", "01010010", "01001010", "01000011", "00111011", "00110100", "00101100", "00100101", "00011101", "00010110", "00001110", "00000111", "00000000" ),
					( "11101111", "11100111", "11011111", "11011000", "11010000", "11001000", "11000000", "10111001", "10110001", "10101001", "10100010", "10011010", "10010010", "10001010", "10000011", "01111011", "01110011", "01101100", "01100100", "01011100", "01010100", "01001101", "01000101", "00111101", "00110110", "00101110", "00100110", "00011110", "00010111", "00001111", "00000111", "00000000" )
				);
					
				data0(2) <= (
					( "00000000", "00000111", "00001111", "00010111", "00011110", "00100110", "00101110", "00110110", "00111101", "01000101", "01001101", "01010100", "01011100", "01100100", "01101100", "01110011", "01111011", "10000011", "10001010", "10010010", "10011010", "10100010", "10101001", "10110001", "10111001", "11000000", "11001000", "11010000", "11011000", "11011111", "11100111", "11101111" ),
					( "00000000", "00000111", "00001110", "00010110", "00011101", "00100101", "00101100", "00110100", "00111011", "01000011", "01001010", "01010010", "01011001", "01100001", "01101000", "01110000", "01110111", "01111111", "10000110", "10001101", "10010101", "10011100", "10100100", "10101011", "10110011", "10111010", "11000010", "11001001", "11010001", "11011000", "11100000", "11100111" ),
					( "00000000", "00000111", "00001110", "00010101", "00011100", "00100100", "00101011", "00110010", "00111001", "01000000", "01001000", "01001111", "01010110", "01011101", "01100101", "01101100", "01110011", "01111010", "10000001", "10001001", "10010000", "10010111", "10011110", "10100110", "10101101", "10110100", "10111011", "11000010", "11001010", "11010001", "11011000", "11011111" ),
					( "00000000", "00000110", "00001101", "00010100", "00011011", "00100010", "00101001", "00110000", "00110111", "00111110", "01000101", "01001100", "01010011", "01011010", "01100001", "01101000", "01101111", "01110110", "01111101", "10000100", "10001011", "10010010", "10011001", "10100000", "10100111", "10101110", "10110101", "10111100", "11000011", "11001010", "11010001", "11011000" ),
					( "00000000", "00000110", "00001101", "00010100", "00011010", "00100001", "00101000", "00101111", "00110101", "00111100", "01000011", "01001001", "01010000", "01010111", "01011110", "01100100", "01101011", "01110010", "01111001", "01111111", "10000110", "10001101", "10010011", "10011010", "10100001", "10101000", "10101110", "10110101", "10111100", "11000010", "11001001", "11010000" ),
					( "00000000", "00000110", "00001100", "00010011", "00011001", "00100000", "00100110", "00101101", "00110011", "00111010", "01000000", "01000111", "01001101", "01010100", "01011010", "01100001", "01100111", "01101110", "01110100", "01111011", "10000001", "10000111", "10001110", "10010100", "10011011", "10100001", "10101000", "10101110", "10110101", "10111011", "11000010", "11001000" ),
					( "00000000", "00000110", "00001100", "00010010", "00011000", "00011111", "00100101", "00101011", "00110001", "00111000", "00111110", "01000100", "01001010", "01010000", "01010111", "01011101", "01100011", "01101001", "01110000", "01110110", "01111100", "10000010", "10001000", "10001111", "10010101", "10011011", "10100001", "10101000", "10101110", "10110100", "10111010", "11000000" ),
					( "00000000", "00000101", "00001011", "00010001", "00010111", "00011101", "00100011", "00101001", "00101111", "00110101", "00111011", "01000001", "01000111", "01001101", "01010011", "01011001", "01011111", "01100101", "01101011", "01110001", "01110111", "01111101", "10000011", "10001001", "10001111", "10010101", "10011011", "10100001", "10100111", "10101101", "10110011", "10111001" ),
					( "00000000", "00000101", "00001011", "00010001", "00010110", "00011100", "00100010", "00101000", "00101101", "00110011", "00111001", "00111111", "01000100", "01001010", "01010000", "01010101", "01011011", "01100001", "01100111", "01101100", "01110010", "01111000", "01111110", "10000011", "10001001", "10001111", "10010100", "10011010", "10100000", "10100110", "10101011", "10110001" ),
					( "00000000", "00000101", "00001010", "00010000", "00010101", "00011011", "00100000", "00100110", "00101011", "00110001", "00110110", "00111100", "01000001", "01000111", "01001100", "01010010", "01010111", "01011101", "01100010", "01101000", "01101101", "01110011", "01111000", "01111110", "10000011", "10001000", "10001110", "10010011", "10011001", "10011110", "10100100", "10101001" ),
					( "00000000", "00000101", "00001010", "00001111", "00010100", "00011010", "00011111", "00100100", "00101001", "00101111", "00110100", "00111001", "00111110", "01000011", "01001001", "01001110", "01010011", "01011000", "01011110", "01100011", "01101000", "01101101", "01110011", "01111000", "01111101", "10000010", "10000111", "10001101", "10010010", "10010111", "10011100", "10100010" ),
					( "00000000", "00000100", "00001001", "00001110", "00010011", "00011000", "00011101", "00100010", "00100111", "00101100", "00110001", "00110110", "00111011", "01000000", "01000101", "01001010", "01001111", "01010100", "01011001", "01011110", "01100011", "01101000", "01101101", "01110010", "01110111", "01111100", "10000001", "10000110", "10001011", "10010000", "10010101", "10011010" ),
					( "00000000", "00000100", "00001001", "00001110", "00010010", "00010111", "00011100", "00100001", "00100101", "00101010", "00101111", "00110100", "00111000", "00111101", "01000010", "01000110", "01001011", "01010000", "01010101", "01011001", "01011110", "01100011", "01101000", "01101100", "01110001", "01110110", "01111011", "01111111", "10000100", "10001001", "10001101", "10010010" ),
					( "00000000", "00000100", "00001000", "00001101", "00010001", "00010110", "00011010", "00011111", "00100011", "00101000", "00101100", "00110001", "00110101", "00111010", "00111110", "01000011", "01000111", "01001100", "01010000", "01010101", "01011001", "01011110", "01100010", "01100111", "01101011", "01110000", "01110100", "01111001", "01111101", "10000001", "10000110", "10001010" ),
					( "00000000", "00000100", "00001000", "00001100", "00010000", "00010101", "00011001", "00011101", "00100001", "00100110", "00101010", "00101110", "00110010", "00110111", "00111011", "00111111", "01000011", "01000111", "01001100", "01010000", "01010100", "01011000", "01011101", "01100001", "01100101", "01101001", "01101110", "01110010", "01110110", "01111010", "01111111", "10000011" ),
					( "00000000", "00000011", "00000111", "00001011", "00001111", "00010011", "00010111", "00011011", "00011111", "00100011", "00100111", "00101011", "00101111", "00110011", "00110111", "00111011", "00111111", "01000011", "01000111", "01001011", "01001111", "01010011", "01010111", "01011011", "01011111", "01100011", "01100111", "01101011", "01101111", "01110011", "01110111", "01111011" ),
					( "00000000", "00000011", "00000111", "00001011", "00001110", "00010010", "00010110", "00011010", "00011101", "00100001", "00100101", "00101001", "00101100", "00110000", "00110100", "00111000", "00111011", "00111111", "01000011", "01000110", "01001010", "01001110", "01010010", "01010101", "01011001", "01011101", "01100001", "01100100", "01101000", "01101100", "01110000", "01110011" ),
					( "00000000", "00000011", "00000110", "00001010", "00001101", "00010001", "00010100", "00011000", "00011011", "00011111", "00100010", "00100110", "00101001", "00101101", "00110000", "00110100", "00110111", "00111011", "00111110", "01000010", "01000101", "01001001", "01001100", "01010000", "01010011", "01010111", "01011010", "01011110", "01100001", "01100101", "01101000", "01101100" ),
					( "00000000", "00000011", "00000110", "00001001", "00001100", "00010000", "00010011", "00010110", "00011001", "00011101", "00100000", "00100011", "00100110", "00101010", "00101101", "00110000", "00110011", "00110111", "00111010", "00111101", "01000000", "01000011", "01000111", "01001010", "01001101", "01010000", "01010100", "01010111", "01011010", "01011101", "01100001", "01100100" ),
					( "00000000", "00000010", "00000101", "00001000", "00001011", "00001110", "00010001", "00010100", "00010111", "00011010", "00011101", "00100000", "00100011", "00100110", "00101001", "00101100", "00101111", "00110010", "00110101", "00111000", "00111011", "00111110", "01000001", "01000100", "01000111", "01001010", "01001101", "01010000", "01010011", "01010110", "01011001", "01011100" ),
					( "00000000", "00000010", "00000101", "00001000", "00001010", "00001101", "00010000", "00010011", "00010101", "00011000", "00011011", "00011110", "00100000", "00100011", "00100110", "00101001", "00101011", "00101110", "00110001", "00110100", "00110110", "00111001", "00111100", "00111111", "01000001", "01000100", "01000111", "01001001", "01001100", "01001111", "01010010", "01010100" ),
					( "00000000", "00000010", "00000100", "00000111", "00001001", "00001100", "00001110", "00010001", "00010011", "00010110", "00011000", "00011011", "00011101", "00100000", "00100010", "00100101", "00100111", "00101010", "00101100", "00101111", "00110001", "00110100", "00110110", "00111001", "00111011", "00111110", "01000000", "01000011", "01000101", "01001000", "01001010", "01001101" ),
					( "00000000", "00000010", "00000100", "00000110", "00001000", "00001011", "00001101", "00001111", "00010001", "00010100", "00010110", "00011000", "00011010", "00011101", "00011111", "00100001", "00100011", "00100110", "00101000", "00101010", "00101100", "00101111", "00110001", "00110011", "00110101", "00111000", "00111010", "00111100", "00111110", "01000000", "01000011", "01000101" ),
					( "00000000", "00000001", "00000011", "00000101", "00000111", "00001001", "00001011", "00001101", "00001111", "00010001", "00010011", "00010101", "00010111", "00011001", "00011011", "00011101", "00011111", "00100001", "00100011", "00100101", "00100111", "00101001", "00101011", "00101101", "00101111", "00110001", "00110011", "00110101", "00110111", "00111001", "00111011", "00111101" ),
					( "00000000", "00000001", "00000011", "00000101", "00000110", "00001000", "00001010", "00001100", "00001101", "00001111", "00010001", "00010011", "00010100", "00010110", "00011000", "00011010", "00011011", "00011101", "00011111", "00100001", "00100010", "00100100", "00100110", "00101000", "00101001", "00101011", "00101101", "00101111", "00110000", "00110010", "00110100", "00110110" ),
					( "00000000", "00000001", "00000010", "00000100", "00000101", "00000111", "00001000", "00001010", "00001011", "00001101", "00001110", "00010000", "00010001", "00010011", "00010100", "00010110", "00010111", "00011001", "00011010", "00011100", "00011101", "00011111", "00100000", "00100010", "00100011", "00100101", "00100110", "00101000", "00101001", "00101011", "00101100", "00101110" ),
					( "00000000", "00000001", "00000010", "00000011", "00000100", "00000110", "00000111", "00001000", "00001001", "00001011", "00001100", "00001101", "00001110", "00010000", "00010001", "00010010", "00010011", "00010101", "00010110", "00010111", "00011000", "00011010", "00011011", "00011100", "00011101", "00011111", "00100000", "00100001", "00100010", "00100100", "00100101", "00100110" ),
					( "00000000", "00000000", "00000001", "00000010", "00000011", "00000100", "00000101", "00000110", "00000111", "00001000", "00001001", "00001010", "00001011", "00001100", "00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111", "00011000", "00011001", "00011010", "00011011", "00011100", "00011101", "00011110" ),
					( "00000000", "00000000", "00000001", "00000010", "00000010", "00000011", "00000100", "00000101", "00000101", "00000110", "00000111", "00001000", "00001000", "00001001", "00001010", "00001011", "00001011", "00001100", "00001101", "00001110", "00001110", "00001111", "00010000", "00010001", "00010001", "00010010", "00010011", "00010100", "00010100", "00010101", "00010110", "00010111" ),
					( "00000000", "00000000", "00000000", "00000001", "00000001", "00000010", "00000010", "00000011", "00000011", "00000100", "00000100", "00000101", "00000101", "00000110", "00000110", "00000111", "00000111", "00001000", "00001000", "00001001", "00001001", "00001010", "00001010", "00001011", "00001011", "00001100", "00001100", "00001101", "00001101", "00001110", "00001110", "00001111" ),
					( "00000000", "00000000", "00000000", "00000000", "00000000", "00000001", "00000001", "00000001", "00000001", "00000010", "00000010", "00000010", "00000010", "00000011", "00000011", "00000011", "00000011", "00000100", "00000100", "00000100", "00000100", "00000101", "00000101", "00000101", "00000101", "00000110", "00000110", "00000110", "00000110", "00000111", "00000111", "00000111" ),
					( "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000" )
				);

	
	Inst_LEDMatrixDriver: LEDMatrixDriver PORT MAP(
		clk => clk,
		sclk => sclk,
		pwm_mode => '1',
		r0 => r0,
		g0 => g0,
		b0 => b0,
		r1 => r1,
		g1 => g1,
		b1 => b1,
		oe => oe,
		latch => latch,
		addr_out => addr_out,
		data => data0,
		rst => rst
	);
	
end Behavioral;

